-- megafunction wizard: %ROM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram

-- ============================================================
-- File Name: digital_rom.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 6.1 Build 201 11/27/2006 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2006 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions
--and other software and tools, and its AMPP partner logic
--functions, and any output files from any of the foregoing
--(including device programming or simulation files), and any
--associated documentation or information are expressly subject
--to the terms and conditions of the Altera Program License
--Subscription Agreement, Altera MegaCore Function License
--Agreement, or other applicable license agreement, including,
--without limitation, that your use is for the sole purpose of
--programming logic devices manufactured by Altera and sold by
--Altera or its authorized distributors.  Please refer to the
--applicable agreement for further details.

LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY digital_rom IS
	PORT (
		address		: IN STD_LOGIC_VECTOR (17 DOWNTO 0);
		clock		: IN STD_LOGIC;
		q		    : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
END digital_rom;


ARCHITECTURE SYN OF digital_rom IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (2 DOWNTO 0);

	COMPONENT altsyncram
        GENERIC (
            clock_enable_input_a		: STRING;
            clock_enable_output_a		: STRING;
            init_file		            : STRING;
            intended_device_family		: STRING;
            lpm_hint		            : STRING;
            lpm_type		            : STRING;
            numwords_a		            : NATURAL;
            operation_mode		        : STRING;
            outdata_aclr_a		        : STRING;
            outdata_reg_a		        : STRING;
            widthad_a		            : NATURAL;
            width_a		                : NATURAL;
            width_byteena_a		        : NATURAL
        );
        PORT (
                clock0	                : IN STD_LOGIC;
                address_a	            : IN STD_LOGIC_VECTOR (17 DOWNTO 0);
                q_a	                    : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
        );
	END COMPONENT;

BEGIN
	q <= sub_wire0(2 DOWNTO 0);

	altsyncram_component : altsyncram
	GENERIC MAP (
		clock_enable_input_a => "BYPASS",
		clock_enable_output_a => "BYPASS",
		init_file => "dig.mif",
		intended_device_family => "Cyclone II",
		lpm_hint => "ENABLE_RUNTIME_MOD=NO",
		lpm_type => "altsyncram",
		numwords_a => 230400,
		operation_mode => "ROM",
		outdata_aclr_a => "NONE",
		outdata_reg_a => "UNREGISTERED",
		widthad_a => 18,
		width_a => 3,
		width_byteena_a => 1
	)
	PORT MAP (
		clock0 => clock,
		address_a => address,
		q_a => sub_wire0
	);

END SYN;
